---------------------------------------------------------------------------------------------------
--
-- Title       : Schematic
-- Design      : design0
-- Author      : Omar Hassan
-- Company     : Lenvo ideapad 5
--
---------------------------------------------------------------------------------------------------
--
-- File        : D:\College\CSE_2_Term_2\Hardware Design\Project\MIPS32-SingleCycle-Processor\design0\design0\compile\Schematic.vhd
-- Generated   : Wed May 15 03:11:24 2024
-- From        : D:\College\CSE_2_Term_2\Hardware Design\Project\MIPS32-SingleCycle-Processor\design0\design0\src\Schematic.bde
-- By          : Bde2Vhdl ver. 2.6
--
---------------------------------------------------------------------------------------------------
--
-- Description : 
--
---------------------------------------------------------------------------------------------------
-- Design unit header --
library IEEE;
use IEEE.std_logic_1164.all;


entity Schematic is 
end Schematic;

architecture Schematic of Schematic is

begin

end Schematic;
